module main;
initial begin
  $display("hello verilog");
  $finish;
end

endmodule
//iverilog hello.v
//vvp a.out